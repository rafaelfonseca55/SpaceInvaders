LIBRARY ieee;
USE ieee.std_logic_1164.all;

Entity COUNTER_UP_DOWN is
Port( CU, CD, RESET, CLK : in std_logic;
		Q : out std_logic_vector(3 downto 0)
        );
End COUNTER_UP_DOWN;

Architecture structure of COUNTER_UP_DOWN is
Component MUX_4 is
Port(A, B : IN STD_LOGIC_VECTOR(3 Downto 0);
        S : In STD_LOGIC;
        Y : Out STD_LOGIC_VECTOR(3 Downto 0));
End Component;

Component ADDER is
Port( A, B : in std_logic_vector(3 downto 0);
        Cin : in std_logic;
        Cout : out std_logic;
        S : out std_logic_vector(3 downto 0)
        );
End Component;

Component REGK is
Port( clk : in std_logic;
		EN : in std_logic;
		D : in std_logic_vector(3 downto 0);
		Q : out std_logic_vector(3 downto 0));
End Component;

signal carry_signal, carry_REG, carry_muxup, carry_muxdown, carry_adder, carry_muxtoadder : std_logic_vector(3 downto 0);

Begin 

U1 : MUX_4 port map (A => "0000", B => "0001", S => CU, Y => carry_muxup);

U2 : MUX_4 port map (A => "0000", B => "1111", S => CD, Y => carry_muxdown);

U3 : MUX_4 port map (A => carry_REG, B => "0000", S => RESET, Y => carry_muxtoadder);

U4 : ADDER port map (A => carry_signal, B => carry_muxtoadder, Cin => '0', S => carry_adder);

U5 : REGK port map (clk => CLK, EN => '1', D => carry_adder, Q => carry_REG);

carry_signal <= carry_muxup or carry_muxdown;

Q <= carry_REG;

End Architecture;

